// Copyright 2018 ETH Zurich and University of Bologna.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.

/*
 // New shifter based on https://github.com/riscv/riscv-bitmanip/blob/main-history/verilog/rvb_shifter/rvb_shifter.v
 *  Copyright (C) 2019  Claire Wolf <claire@symbioticeda.com>
 *
 *  Permission to use, copy, modify, and/or distribute this software for any
 *  purpose with or without fee is hereby granted, provided that the above
 *  copyright notice and this permission notice appear in all copies.
 *
 *  THE SOFTWARE IS PROVIDED "AS IS" AND THE AUTHOR DISCLAIMS ALL WARRANTIES
 *  WITH REGARD TO THIS SOFTWARE INCLUDING ALL IMPLIED WARRANTIES OF
 *  MERCHANTABILITY AND FITNESS. IN NO EVENT SHALL THE AUTHOR BE LIABLE FOR
 *  ANY SPECIAL, DIRECT, INDIRECT, OR CONSEQUENTIAL DAMAGES OR ANY DAMAGES
 *  WHATSOEVER RESULTING FROM LOSS OF USE, DATA OR PROFITS, WHETHER IN AN
 *  ACTION OF CONTRACT, NEGLIGENCE OR OTHER TORTIOUS ACTION, ARISING OUT OF
 *  OR IN CONNECTION WITH THE USE OR PERFORMANCE OF THIS SOFTWARE.
 *
*/

////////////////////////////////////////////////////////////////////////////////
// Engineer:       Matthias Baer - baermatt@student.ethz.ch                   //
//                                                                            //
// Additional contributions by:                                               //
//                 Igor Loi - igor.loi@unibo.it                               //
//                 Andreas Traber - atraber@student.ethz.ch                   //
//                 Michael Gautschi - gautschi@iis.ee.ethz.ch                 //
//                 Davide Schiavone - pschiavo@iis.ee.ethz.ch                 //
//                 Halfdan Bechmann - halfdan.bechmann@silabs.com             //
//                                                                            //
// Design Name:    ALU                                                        //
// Project Name:   RI5CY                                                      //
// Language:       SystemVerilog                                              //
//                                                                            //
// Description:    Arithmetic logic unit of the pipelined processor           //
//                                                                            //
////////////////////////////////////////////////////////////////////////////////


module cv32e40x_alu import cv32e40x_pkg::*;
(
  input  logic              clk,
  input  logic              rst_n,
  input  alu_opcode_e       operator_i,
  input  alu_shifter_t      shifter_i,
  input  logic [31:0]       operand_a_i,
  input  logic [31:0]       operand_b_i,

  output logic [31:0]       result_o,
  output logic              comparison_result_o,

  // Divider interface towards CLZ
  input logic               div_clz_en_i,
  input logic [31:0]        div_clz_data_i,
  output logic [5:0]        div_clz_result_o,

  // Divider interface towards shifter
  input logic               div_shift_en_i,
  input logic [5:0]         div_shift_amt_i,
  output logic [31:0]       div_op_a_shifted_o
);

  //logic [31:0] operand_a_rev;
  
  // bit reverse operand_a for left shifts and bit counting
 /* generate
    genvar k;
    for(k = 0; k < 32; k++)
    begin : gen_operand_a_rev
      assign operand_a_rev[k] = operand_a_i[31-k];
    end
  endgenerate
*/
  logic [31:0] operand_b_neg;

  assign operand_b_neg = ~operand_b_i;


 ////////////////////////////////////////
  //  ____  _   _ ___ _____ _____       //
  // / ___|| | | |_ _|  ___|_   _|      //
  // \___ \| |_| || || |_    | |        //
  //  ___) |  _  || ||  _|   | |        //
  // |____/|_| |_|___|_|     |_|        //
  //                                    //
  ////////////////////////////////////////

  logic        shifter_rotate;
  logic        shifter_rshift;
  logic        shifter_arithmetic;
  logic        shifter_operand_tieoff; // Ties shifter oprand a to 1 and b to 0. Used for some single bit operations.

  logic [31:0] shifter_bext_result;
  logic [31:0] shifter_bset_result;
  logic [31:0] shifter_bclr_result;
  logic [31:0] shifter_binv_result;

  logic [63:0] shifter_tmp;
  logic [5:0]  shifter_shamt;  // Shift amount
  logic [31:0] shifter_result; // Shift right
  logic [31:0] shifter_aa, shifter_bb;


  assign shifter_rotate         = (div_shift_en_i) ? 1'b0 : shifter_i.rotate;
  assign shifter_rshift         = (div_shift_en_i) ? 1'b0 : shifter_i.rshift;
  assign shifter_arithmetic     = (div_shift_en_i) ? 1'b0 : shifter_i.arithmetic;
  assign shifter_operand_tieoff = (div_shift_en_i) ? 1'b0 : shifter_i.operand_tieoff;


  assign div_op_a_shifted_o = shifter_result;
  always_comb begin
    //Can mess up the divider?
    shifter_shamt = div_shift_en_i ? {1'b0, div_shift_amt_i[4:0]} : {1'b0, operand_b_i[4:0]};
    shifter_aa = (shifter_operand_tieoff) ? 32'h1 : operand_a_i;

    //TODO: might not be nessessary, ask what shifter_operand_tieoff does!
    //For the moment make sure we set correct shifter_aa value:
    //if ((operator_i == ALU_B_SH1ADD) || (operator_i == ALU_B_SH2ADD) || (operator_i == ALU_B_SH3ADD)) shifter_aa = operand_a_i; //Try to take this out!

    //OBSOBS!
    
    if (shifter_rshift) begin
      // Treat right shifts as left shifts with corrected shift amount
      shifter_shamt = -shifter_shamt;
    end

    //In case of a SHxADD operation set shifter_shamt accordingly
   // if (operator_i == ALU_B_SH1ADD && !div_shift_en_i) shifter_shamt =  $unsigned(1);
   // if (operator_i == ALU_B_SH2ADD && !div_shift_en_i) shifter_shamt =  $unsigned(2);
   // if (operator_i == ALU_B_SH3ADD && !div_shift_en_i) shifter_shamt =  $unsigned(3);
    
    
    if (shifter_operand_tieoff) begin
      shifter_bb = 32'h0;
    end else if (shifter_arithmetic) begin
      shifter_bb = shifter_rotate ? operand_a_i : {32{operand_a_i[31]}};
    end else begin
      shifter_bb = shifter_rotate ?          '1 : '0;
    end

  end

  always_comb begin
    shifter_tmp = {shifter_bb, shifter_aa};
    shifter_tmp = shifter_shamt[5] ? {shifter_tmp[31:0], shifter_tmp[63:32]} : shifter_tmp;
    shifter_tmp = shifter_shamt[4] ? {shifter_tmp[47:0], shifter_tmp[63:48]} : shifter_tmp;
    shifter_tmp = shifter_shamt[3] ? {shifter_tmp[55:0], shifter_tmp[63:56]} : shifter_tmp;
    shifter_tmp = shifter_shamt[2] ? {shifter_tmp[59:0], shifter_tmp[63:60]} : shifter_tmp;
    shifter_tmp = shifter_shamt[1] ? {shifter_tmp[61:0], shifter_tmp[63:62]} : shifter_tmp;
    shifter_tmp = shifter_shamt[0] ? {shifter_tmp[62:0], shifter_tmp[63:63]} : shifter_tmp;
  end

  assign shifter_result      = shifter_tmp[31:0];

  assign shifter_bext_result =       32'h1 &  shifter_result;
  assign shifter_bset_result = operand_a_i |  shifter_result;
  assign shifter_bclr_result = operand_a_i & ~shifter_result;
  assign shifter_binv_result = operand_a_i ^  shifter_result;


  //////////////////////////////////////////////////////////////////////////////////////////
  //   ____            _   _ _   _                      _      _       _     _            //
  //  |  _ \ __ _ _ __| |_(_) |_(_) ___  _ __   ___  __| |    / \   __| | __| | ___ _ __  //
  //  | |_) / _` | '__| __| | __| |/ _ \| '_ \ / _ \/ _` |   / _ \ / _` |/ _` |/ _ \ '__| //
  //  |  __/ (_| | |  | |_| | |_| | (_) | | | |  __/ (_| |  / ___ \ (_| | (_| |  __/ |    //
  //  |_|   \__,_|_|   \__|_|\__|_|\___/|_| |_|\___|\__,_| /_/   \_\__,_|\__,_|\___|_|    //
  //                                                                                      //
  //////////////////////////////////////////////////////////////////////////////////////////

  logic        adder_op_b_negate;
  logic [31:0] adder_op_a, adder_op_b;
  logic [32:0] adder_in_a, adder_in_b;
  logic [31:0] adder_result;
  logic [33:0] adder_result_expanded;

  assign adder_op_b_negate = (operator_i == ALU_SUB);

  // prepare operand a
  assign adder_op_a = operand_a_i;  //(operator_i == ALU_ADD || operator_i == ALU_SUB) ? operand_a_i : shifter_result;

  // prepare operand b
  assign adder_op_b = adder_op_b_negate ? operand_b_neg : operand_b_i;

  // prepare carry
  assign adder_in_a = {adder_op_a, 1'b1};
  assign adder_in_b = {adder_op_b, adder_op_b_negate};

  // actual adder
  assign adder_result_expanded = $unsigned(adder_in_a) + $unsigned(adder_in_b);
  assign adder_result = adder_result_expanded[32:1];

  
  //////////////////////////////////////////////////////////////////
  //   ____ ___  __  __ ____   _    ____  ___ ____   ___  _   _   //
  //  / ___/ _ \|  \/  |  _ \ / \  |  _ \|_ _/ ___| / _ \| \ | |  //
  // | |  | | | | |\/| | |_) / _ \ | |_) || |\___ \| | | |  \| |  //
  // | |__| |_| | |  | |  __/ ___ \|  _ < | | ___) | |_| | |\  | and min/max  //
  //  \____\___/|_|  |_|_| /_/   \_\_| \_\___|____/ \___/|_| \_|  //
  //                                                              //
  //////////////////////////////////////////////////////////////////

  logic is_equal;
  logic is_greater;     // handles both signed and unsigned forms
  logic cmp_signed;

  assign cmp_signed = (operator_i == ALU_GES) || (operator_i == ALU_LTS) || (operator_i == ALU_SLTS) || (operator_i == ALU_B_MIN) || (operator_i == ALU_B_MAX);
  assign is_equal = (operand_a_i == operand_b_i);
  assign is_greater = $signed({operand_a_i[31] & cmp_signed, operand_a_i}) > $signed({operand_b_i[31] & cmp_signed, operand_b_i});

  // generate comparison result
  logic cmp_result;

  always_comb
  begin
    cmp_result = is_equal;
    unique case (operator_i)
      ALU_EQ:            cmp_result = is_equal;
      ALU_NE:            cmp_result = ~is_equal;
      ALU_GES, ALU_GEU:  cmp_result = is_greater | is_equal;
      ALU_LTS, ALU_SLTS,
      ALU_LTU, ALU_SLTU: cmp_result = ~(is_greater | is_equal);

      default: ;
    endcase
  end

  assign comparison_result_o = cmp_result;

  // generate min/minu and max/maxu result:
  logic [31:0] min_minu_result;
  logic [31:0] max_maxu_result;

  assign min_minu_result = (!is_greater) ? operand_a_i : operand_b_i;
  assign max_maxu_result = (is_greater) ? operand_a_i : operand_b_i;

 
  /////////////////////////////////////////////////////////////////////
  //   ____  _ _      ____                  _      ___               //
  //  | __ )(_) |_   / ___|___  _   _ _ __ | |_   / _ \ _ __  ___    //
  //  |  _ \| | __| | |   / _ \| | | | '_ \| __| | | | | '_ \/ __|   //
  //  | |_) | | |_  | |__| (_) | |_| | | | | |_  | |_| | |_) \__ \_  //
  //  |____/|_|\__|  \____\___/ \__,_|_| |_|\__|  \___/| .__/|___(_) //
  //                                                   |_|           //
  /////////////////////////////////////////////////////////////////////

  logic [31:0] div_clz_data_rev;
  logic [31:0] clz_data_in;
  logic [4:0]  ff1_result; // holds the index of the first '1'
  logic        ff_no_one;  // if no ones are found
  logic [ 5:0] cpop_result_o;
  //logic [31:0]  clmul_result;

  assign clz_data_in = (operator_i == ALU_B_CTZ) ?  div_clz_data_rev : div_clz_data_i;

  generate
    genvar l;
    for(l = 0; l < 32; l++)
    begin : gen_div_clz_data_rev
      assign div_clz_data_rev[l] = div_clz_data_i[31-l];
    end
  endgenerate

  cv32e40x_ff_one ff_one_i
  (
    .in_i        ( clz_data_in ),
    .first_one_o ( ff1_result ),
    .no_ones_o   ( ff_no_one  )
  );

  // Divider assumes CLZ returning 32 when there are no zeros (as per CLZ spec)
  assign div_clz_result_o = ff_no_one ? 6'd32 : ff1_result;
 

  // CPOP
  cv32e40x_alu_b_cpop alu_b_cpop_i
    (.operand_i (operand_a_i),
     .result_o  (cpop_result_o));

  /////////////////////////////////
  //  carryless multiplication   //
  /////////////////////////////////
//ADDED - FRAME CLMUL/H/R version framework
  /*
  logic [31:0] operand_a_rev;
  logic [31:0] operand_b_rev;
  
  logic [31:0] operand_a_clmul;
  logic [31:0] operand_b_clmul;
  
  logic [31:0] clmul;
  logic [31:0] clmulr;
  logic [31:0] clmulh;
  
  for (genvar k = 0; k < 32; k++) begin
    assign operand_a_rev[k] = operand_a_i[31-k];
    assign operand_b_rev[k] = operand_b_i[31-k];
  end

  assign operand_a_clmul = (operator_i != 2'b00) ? operand_a_rev : operand_a_i;
  assign operand_b_clmul = (operator_i != 2'b00) ? operand_b_rev : operand_b_i;

  for (genvar k = 0; k < 32; k++) begin
    assign clmulr[k] = clmul[31-k];
  end

  assign clmulh = {1'b0, clmulr[31:1]};
  */
//ADDED framework - FINISHED  

  //ADDED YouTube different result
  logic [1:0] operator_clmul;
  logic [31:0] clmul_result;

  assign operator_clmul = (operator_i == ALU_B_CLMUL) ? 2'b00 : (operator_i == ALU_B_CLMULH) ? 2'b01 : 2'b10;
  
  //ADDED Youtube different result finished
  cv32e40x_alu_b_clmul alu_b_clmul_i
    (.op_a_i (operand_a_i),
     .op_b_i (operand_b_i),
     .operator_i(operator_clmul),
     .result_o  (clmul_result)
    // .result_o(clmul)
      );

  /*
  /////////////////////////////////
  //    min/max instructions     //
  /////////////////////////////////
  logic [31:0]  min_result;
  logic [31:0]  minu_result;
  logic [31:0]  max_result;
  logic [31:0]  maxu_result;
  assign min_result  = (  $signed(operand_a_i) <   $signed(operand_b_i)) ? operand_a_i : operand_b_i;
  assign minu_result = ($unsigned(operand_a_i) < $unsigned(operand_b_i)) ? operand_a_i : operand_b_i;
  assign max_result  = (  $signed(operand_a_i) >   $signed(operand_b_i)) ? operand_a_i : operand_b_i;
  assign maxu_result = ($unsigned(operand_a_i) > $unsigned(operand_b_i)) ? operand_a_i : operand_b_i;
*/

////////////////
// shift add  //
////////////////

  logic [31:0] shXAdd;
  logic [31:0] shX;
  
  assign shX = (operator_i == ALU_B_SH1ADD) ? operand_a_i << 1 : (operator_i == ALU_B_SH2ADD) ? operand_a_i << 2 : operand_a_i << 3; 
  
  assign shXAdd = shX + operand_b_i;
 
  
  ////////////////////////////////////////////////////////
  //   ____                 _ _     __  __              //
  //  |  _ \ ___  ___ _   _| | |_  |  \/  |_   ___  __  //
  //  | |_) / _ \/ __| | | | | __| | |\/| | | | \ \/ /  //
  //  |  _ <  __/\__ \ |_| | | |_  | |  | | |_| |>  <   //
  //  |_| \_\___||___/\__,_|_|\__| |_|  |_|\__,_/_/\_\  //
  //                                                    //
  ////////////////////////////////////////////////////////

  always_comb
  begin
    result_o   = '0;

    unique case (operator_i)
      // Standard Operations
      ALU_AND:  result_o = operand_a_i & operand_b_i;
      ALU_OR:   result_o = operand_a_i | operand_b_i;
      ALU_XOR:  result_o = operand_a_i ^ operand_b_i;

      // Adder Operations
      ALU_ADD,
      ALU_SUB : result_o = adder_result;

      // Shift Operations
      ALU_SLL,
        ALU_SRL, ALU_SRA:  result_o    = shifter_result;

      // Non-vector comparisons
      ALU_SLTS,  ALU_SLTU: result_o    = {31'b0, comparison_result_o};

      // RV32B Zca instructions
      // TODO:OE: Investigate sharing ALU adder and shifter
    
       //SOMETHINGS!!!
      ALU_B_SH1ADD, ALU_B_SH2ADD, ALU_B_SH3ADD: result_o = shXAdd;  //adder_result; //shifter_result;
      //ALU_B_SH1ADD: result_o = (operand_a_i << 1) + operand_b_i;
      //ALU_B_SH2ADD: result_o = (operand_a_i << 2) + operand_b_i;
      //ALU_B_SH3ADD: result_o = (operand_a_i << 3) + operand_b_i;


      // Zbb
      ALU_B_CLZ, ALU_B_CTZ: result_o   = {26'h0, div_clz_result_o};
      ALU_B_CPOP:           result_o   = {26'h0, cpop_result_o};
      
      ALU_B_MIN, ALU_B_MINU:  result_o = min_minu_result;
      ALU_B_MAX, ALU_B_MAXU:  result_o = max_maxu_result;
     
      ALU_B_ANDN:           result_o   = operand_a_i & ~operand_b_i;
      ALU_B_ORN:            result_o   = operand_a_i | ~operand_b_i;
      ALU_B_XNOR:           result_o   = operand_a_i ^ ~operand_b_i;

      ALU_B_ORC_B:          result_o   = {{(8){|operand_a_i[31:24]}},
                                        {(8){|operand_a_i[23:16]}},
                                        {(8){|operand_a_i[15:8]}},
                                        {(8){|operand_a_i[7:0]}}};

      ALU_B_REV8:           result_o = {operand_a_i[7:0],
                                        operand_a_i[15:8],
                                        operand_a_i[23:16],
                                        operand_a_i[31:24]};
      ALU_B_ROL,
        ALU_B_ROR:            result_o = shifter_result;

      ALU_B_SEXT_B:         result_o   = {{(24){operand_a_i[ 7]}}, operand_a_i[ 7:0]};
      ALU_B_SEXT_H:         result_o   = {{(16){operand_a_i[15]}}, operand_a_i[15:0]};

      // Zbs
      ALU_B_BSET:           result_o   = shifter_bset_result;
      ALU_B_BCLR:           result_o   = shifter_bclr_result;
      ALU_B_BINV:           result_o   = shifter_binv_result;
      ALU_B_BEXT:           result_o   = shifter_bext_result;

      // Zbc
      ALU_B_CLMUL, //:           result_o  = clmul;
      ALU_B_CLMULH, //:          result_o  = clmulh;
      ALU_B_CLMULR:          result_o  = clmul_result;  //clmulr;
      
      

      default: ; // default case to suppress unique warning
    endcase
  end

endmodule // cv32e40x_alu
